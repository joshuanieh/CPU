module Control(
    Op_i,
    ALUOp_o,
    ALUSrc_o,
    RegWrite_o
);

